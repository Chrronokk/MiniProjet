antoine@localhost.8050:1513084798