xph2sei409@cimeld11.2808:1523962287