antoine@localhost.21783:1513084798