xph2sei409@cimeld11.24773:1523962287