xph2sei409@cimeld11.15611:1523962287