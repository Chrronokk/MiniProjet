library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package programme is

  type B32 is array (0 to 51) of std_logic_vector(7 downto 0);  -- mémoire interne

  constant prog : B32 :=
    ("00000000","00000000","00000000","00000000",
     "11111111","11111001","00001000","00010011",  --ADDI r20,111111111111->r16
     "00000000","00010000","10000000","10010011",  --ADDI r1,1->r1
     "00000001","00000000","10100000","00100011",  --SW r16,mem(r1)
     "00000000","00000000","10000010","00000011",  --LB mem(r1),r4
     "00000000","00000000","11000010","10000011",  --LBU mem(r1),r5
     "00000000","00000000","10010011","00000011",  --LH mem(r1),r6
     "00000000","00000000","11010011","10000011",  --LHU mem(r1),r7
     "00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000");

  
  

end programme;
