antoine@localhost.29405:1513084798