xph2sei409@cimeld11.15820:1523962287