xph2sei409@cimeld11.2787:1523962287