library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package programme is

  type B32 is array (0 to 67) of std_logic_vector(7 downto 0);  -- mémoire interne

  constant prog : B32 :=




    ("00000000", "00000000", "00000000", "00000000",
     "00000000", "01110000", "00000101", "00010011",  --ADDI 111 -> r10
     "00000000", "01000000", "00000100", "10010011",  --ADDI 100 -> r9
     "00000000", "10100100", "10100001", "00100011",  --SW r10 -> mem(r9)+2
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "00100100", "10101000", "00000011",  --LW mem(r9)+2 -> r16
     "00000100", "00011000", "01100110", "00010011",  --ORI r16,1000001 -> r20
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "10001010", "00000010", "01100111",  --JALR:(PC<-R0+10)&(R4<-PC+4)     ,
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "00000000", "00000000", "00000000",
     "00000000", "00000000", "00000000", "00000000");




end programme;
